0
1
(1;1.28941) = (2;1.7853)

